��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��6�L�h�p@�
�D�i�����[�B$�N-ɛ#R \h��/6)��nJ�z)g~�HZE�x��{R6���-���r���)n�vl�ɒ-�)E��ww85��� ��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O����w��=�3�n����0:��q�q��%�J�`���l�d6��p�y~ �z8`���K�<��I��ؕ���~�aVw���}Ẃ���:j6\�(o%5��Y�~%$]���ZGfa�XC7�b@�t	aJ�:�?�WG���#�W��\j@ϝ+�'}V�5j���AVЪv_O.&�4v�Er��z�=�4"�c\s��J>��m_��^,�2A��S5���	(hN�X������=4�Cg��Uf9���jɫF�[��`�Wu�Ͷ+��AEM|�W��]�L�[y�ɺW���c�Xn�W�afW�*OH���r_�Q�ut�iߎi*��{��bϢP\͏���:�ޓٗ� �qs�n�һ(HR���wI��ܙ�wi��|;���������`��cCĞ�$S�h��@QI�
n&�]��3rm}r.vX�դ�W��]b�s�v,�Z"�� a�O���G��B��e��n���+Δ}183ge��I���l_�e��&~����⎅��'�̳~�z)����[S�v��	1+��	Bb0�J���}���1
��̸}E)�'��t�^c'ߓ�%�<�Ek8?H�5��2kp��Xe��& Q��m0U�E��w�g�d8g�?c����cB	�VE�<ӽ���p'��l������q.�����ʂ�#��<�S�6����[+��#\�^��ț�����`�X-������M����yQV�uY���z��S�8gc�匾vtޓ���23�B�t���1�C&B:���O�r�	8�����d^dƌN,b�.0c�׻:5 �L�$2H�����C�A��#��;�!��/&oL2�B��/�Ra��9��g2�AU�Մ���5�I���%[D��-�I�˶@'#ضc�����_H&[�I8�^��R��Y�ֱʋ�O^��~N�߽^菇ܪ�����t��t�9/���T������m�$w��6ӑ̮�W��� �Y�9
���
����
��1���M��S���5��qt���H'؇�
6���/��E��s��-߾8qG~�L #�a:���Y.�=p%�
�c�?)q�gc{�BP�ݹ,����y^FZL��f�\)lN���L�$IK tn���G���0�L�����Nɷy>D)�F!��(uE͍� ���GT!�s8��������)�V��,w�^�3�w� MpU�ɇW���j�,���yƝ6�n0��k�'sC�ڟyn�mj��<����W�.A���ߎ<���\`�xW������A�%�T*o�#�2�u�5rJ1tUG�a����Dʊͅ>�3�.���5��e�Q��yP�u��u�����٭�B��u^ԭtgp�K���\�>���<���/Y�2�7d�D�p����s5��$C�?Q~�I��~�H0�0���DI�ܼR���%��v` U�}��в�3��1%��AS԰&�H\���=8@��P߳�,N�'�'g�~+�Cd'i&�.����[8o�E�?�W�M\I�����.@�=A�O�;�mP_�-Ꮇ��I�k�G�飺�S�ug��],�P^�t<2�s�Q�=�1� Q�er't#�#�QT�T�}����ʡ��f�:kc��'�N����5���|'����Gq`�%�`��s��E�9�9o<��Ĩ_W��l8d@��Pȋ�9D��ʄ��OR�LLN�V�@v�@}�_��z����e�a<L��3�ޱcŽH�u�?-�k�����c�?����ι�Ot$sKĉ�)1!M���SMvy�Y+��Lj}T�>Y��U]�r���F��hy�U�x�gn���x볮��b�����[���%�s
�����S�#,2HK1i�D�.�N��U�ӢAv$9��ϠJ��������x�6�dΎy}���V��,/�[t�BiP
7D>
��k��R(��C�����s�b�`��r��)2�r'.��k, ���@�n��*�+���+@��ו��� 
�Ų����}t��� ;f��M�	��,U��K��̼�+��.��=�ț\�S0Q���"j��RE���Qt-�`-Ak��=�W�Za�u��r.�͘�ŉciZ��(� l	`'.E%�W�1��)����1���V�l<����h�`d��K�v��kz�FaX�0�ä���YЬ��3_{k�T��կ�L@;���2M�*��`5�,;�C�x�3�%�m��6��Zkyl1���!J�4A�P�9��O�ux^���\k�>���c���*� ��1-#Rެ:=�]v@o�(jgE�R���|�rJ��Pl��C����Er�zq�2�G�
[��v�gb�F���ߜs �L��Y7�s�,�2z􌸵L{s�|�]����q�� ��atn+�w�0ZD�ʒo�R�A�c��p��F�>A�t���W��*|�Ό�8�wcB��=�i�ùȕ�p���{p\_)��%��E�$T��3)���	��:t:���,��_ �X�&=�>�׾�+���3Ax_u���2��Z2�FFCNLQ� p5�g��K�U&�r0�f��ž9'��- �U5��5$RN�:to/��H�!�����B����I�Ir\�z���AA��s����Tp�.�a�B�7S�"�����xy�
��t�8�uX,�3���H;w=+O��J�/�:�OUKR�M���<K��b��o7��^�d@�;�j�J�:]}B�G1�����\�<}�)�p¦��4�w���n{ǣ�D�S)tг:�M2Dz�v�Ϋ����W�W�Sa�N��Z�����j7�%�p���A�|���ZX֘lk0,� O"~F�A����E�l������2��s�#��^��0�C��ў\2K=����"��SvP�H��;�fTF,�(��!$���Z,:!�{qe��lh,hR� °��$W:1��M$�>��Q�*��;,.�C���1�O"m�P����R(��5=̜��՗�1/��z��

*���)lF���������ϺĂR|1?��i�bz�9]��{����җ��ߧa�\�_�:��q���C}�e��I�7fj ��i
�C��xO�+Ȋ
dpNe����j��R�: �N��H\w�q��4wl!�vJ'jd=�����.�ۛ�{�|x޸kCR4[j�:v��5�k���n�������UM����&Q���a����GZ���d��ڴ5��l�| gJ��������k��U��׀�v)^��I��!�62 ��Q\�v���8)�B���0O@��z<��%LY=}�h+4�@���l "ou�;�H�7�
A���K�)��2�碋���}']�����r��8q�+y��ǁ��x�+=
��y���~Ɛ���K�+A�`υ2�ם�w1E7�9��u��~#����]X;�s���W|�1���x}�t���6�h-�%�(����������Q&�"�:��aM��9d劑Et%��*
L|�;���k0E0?�Э�k�aL%����3!8Y�1�}^��5q�ɴ�pN꧰�ꆽ���-�m�ߡǋ��%��V���j�m[QxK����{ +p'iI^��k}��9~S�Ϲ�+��2�^Mf����r���`���t�̕��Y����{�502�����!`Am���o� ��}��{��m翏����ŀ^�O~����;�ke���}����_;T���jU"H����D�{3�E^^���HFk�";�%�(1����ay�L�K��U����*w��/��9_"��ϨS�*��V�P����(������ۢ�[�Db���Ԛ��@`�wɚ��2�;���u�%:S�
����ko�ǟUŞ叏4;��^ү�e��!��ք�rik�Z&(³l��wktu���hU"�p�ْ����w����cƸ7�]{�� N���o+S��z]J����~W��� K���v&6������/�㛙�\w�1����|�xe45>2�B$��5��
��3풯� ��b�q�9��J]<ms7Q�(���%�I�H÷�T�-ޞ���&�Q� �������қ�=��w�g�V�)��C����q�*�P�~1t�[���Ap߬%�p�Dv';�bMy��hT��P��E���}{O�zՈ�j�w�<��#4���ΉQD+J��&]Q��[m���q�M3�ʂ�t�d�L�u����=D���!�hŽ8S����ݿ٢�\D1�������!dE�w��%:/Q;~���R�AQ>n�E������؆1�ᛸ�6����Ls�0����=�E%�ƶ�(W�2�CMt�$z���=�ٟ�gXi����H;|���m��P"�O8f.���[J�pY[AlK{��栣A���["�a^YG��KqZ�1Xe�.�)?1ɹ��[zm��H2(Q:7o2�O�;�G��2�\��\R�C0	�X(~�t�<��zf�*?��Ͻ���vt���l���P;� #b��!���5~�[;P�|�AX���+/b�e_eB����R��r�3��!��Q^q:�pg	N����c�de���S�cB�Lܦ�߂K֍�/A��r����0	�)�\Vg����l�� drO�D��v;���凋Q{��i��!���5�`G� ?V&J;]�� �	&�92�Y�K)��4�Ĥ�4Q���$�x�M~Ÿ�ٔ���2y��8	o��Dx|f�r�fC�\8�1��n�SQi�9��vF$;��H> 5# �Y�|��V��md���;������z��8����+{;��S�����ǰd���֭�H� ���Uv�*il���l�9�ݹG�lZJ��"�n}�l��z���K�ƽ?����m��s$�鋡��mQ��k�T��zz|rL�i w`�%�/,E(a�N-��Y(`����������K�U������ ~=1��F~�q/�t���n#!��a#���͹Uȅ�����2 (�[�I�9/�Y���w���������qT�Ɉ�|��8�@���C{�$9hD���iu5� �X��x�wvF��`(#0�!�
�Vo�VJ��U0a�o.RҢ��a�t
,H訹�U�x��'� dP�{k�?H��B<�k���cE'�{?b	/X>�圑���Wli�`ь!���i�]���q�[�Q�>͐���L.5=�:
:ss�6�G��8v�T؄����2���҃�Ys`Ǟ3�ᶣ?~Iy�<�	1vol��p�&4&;�+��^���*	�f�|o�g{�Mݩ�o������-�f�[�*4Dz�Lhi���Q	�-�y�(�