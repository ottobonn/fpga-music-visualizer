��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��6�L�h�p@�
�D�i�����[�B$�N-ɛ#R \h��/6)��nJ�z)g~�HZE�x��{R6���-���r���)n�vl�ɒ-�)E��ww85��� ��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O����w��=�3�n��Ht�#w!{��4�6��QKv�c�0F}ͣ�
��u��-F���������V��|�80 ���O�IG�r��� �:�@���{���ӾZ����\Ƌ�ב�,��{�Y�c�i|$g*R�7�����
��M����q���
n�6& �ϝ�s/��b�ԥasV��0�� �P��/{!G6��F�5���
q�!Y�
8�%F�w�P��vx�M�Ju�&G��|K��M��N��� �r��n.Z7I\���I������	d��6��Q	'���6(QEw��"�_�^���U.�i�d8�`����tBB  �cn�j{�`A�:t҃;/�jƵ�k���xV:ܰ�N��E�.�L���
��]�����tZ�o���=Y����� H=&��g�(��#(�R��~��j7�[����/C��k�o8�i��c���Ճ�Z'ޫ�YS��#^{SM	`�x���>�T=(q���<���
�'�y"n��	җ;)1�ؑ+y�촐L�E���x�^%���NN�ś����$��к,IM)�4q����5�!�œi(*~��<����!^���z=!�k�����0���.`�({��K�և��	��R{�&����Hny�o5��9y���(}��QwS��@յ����J�j&l�B�5�_wl4�y�1.=ǃ�6Ҽ i���{�|�Z�0�"���_c���;�O3f��P����I�WM��,Tq�d-�>FC��̅	�^ ���*ȧҖӀ��=�[%��#~G䱁�}N��^�i�9x��8���VR��vM!)�;�;�4��"|;1���I~���	����0`����@d\E��h?�ƼI�	��%zJ�*C~�@��ѷ�Kc=�]�	�I��s�����S��m\%U ��� �م�h!�&�U$�dԺ��v���$�����bl�Z�jUn���R.��lڰ�*�g��%��f���Q-�Ja����~��Н�=����K��W�a����`Z���6�-��, |��}M�*����6/h�t�{�ۑd�/+��m�����n}*�X��9�,��h(š"]D.c�'B$�@&Ў�3��p89�?Io��J9U�6�˃=0�5�&[��-�q<~��,���7����
�-�h~�+IL�5�}��9��:^[��<=J�^%M���d��9_�SL ~:[��O�dY%.����:Tˆ&��Qy��[F�4I��Q���w�CfR�֧������z�h��o)N��?���K�HgX�� g\Ƈ7�mL�����ڭ���>L̠���0h�` �P�,Lܖ���F�Wd4&�h��@�_&���<ΙX&۞��������7�{���-��NQ�����H��q���R,�ct$
�Ǽ_��(_���?d_���6LZE��X�JM ���
�-�n�� ��(8f�Ѷ�Ύ�^��G*����9,�\����_?�<����)��%��ka����$E�&���d�,o�p�d.��d�KY�D���0��It�<������lW5gE(>:
�������� ���R(��Tr�-&�B4P_jW��|cZX����):Zxȿ"J�b8Ԇ�F��Q�����G�6���Mſ��m`�x��C�l�-h�)@z�Օ%(�\j#�����B�G�.u3�%Q"$t�������igm1OB^~.�������w=�
�9&�A��k;J�cH�������s|��Փ/��ó� ݀��>��ZB����浗x�I�F�M��Va����,��ɦ0�JL�Ae^�a�l
7�e��Y�G1�/-"#���Զ)��5��X��(����G�y]��ρ�����-��Enk��BiUYf*��^�r��,��ǎ[.�ܧ���������?�2���N�1�8�"0=�oT֮]�q݁ n2�R��h�����x���I;��([�H�JG��[ZK���������U��L?kE����F`����kT`af.��Hg0T`����/����ص�1D�m������Yϖd��'Z9{`���>�5�����ӣ��Uݯ8x�>؆��}z�P����S��o��t�
<^���{&vEq�"����$1�]�F�^f��)��"Z��:rh����3I��yK�V6t@^�������S���W���}p8�h�1������d��m�0(�m~�l!B�Q�䭎�w��(E���ֺ�ō�-��q�!���a%����9������U��n02���G�k�6X֭)��~{�ϑH��`�~���:��짰�mt�KK|so7�r���V���������(�"Y$�$�	��/��赎*k�C���̊$����j�)�>Kҽ�m���/�*�b�~�4z�4K�R^'?��\a\j�$������7^�=؊rw�\�@�Ct��yX��/L�-x�XZ�ے"g�gǩ����_S`t��=��_�>�1K��'���jl#K$�^��ÁmK!R��ݷ�->u:��9����݇X̑�ܞ�3�v�G��zH��Q~�vw�~���8�L����N �˒:3櫘���+@1w���7��<cE��x���Ϭ���{�?��?�s�″f�0_QO����οbp��I��[oEo;�������1�yG� I`���Lx~r�Z�sM:�J�K�����|���Δ�]��Bo皝�ER���s>�|�;�2ϿˀzZ�������lh����	�������8s�[�}X��v�m�`�X
�?��ӂ�����I ��B,-��<<� ��f$��@^�d/IA�$���բ0 ��kS�o=�I���`^���Zy�(�e�v���%�N�y��V�/�xa��Z2�P�>�5�i�q�Ė�K	Ȇ������[�[�� ¿͂�+$0�˩������>� l�+|��,������J���bЀ�.}���G�zQ���${��LG�B#�֨3/�e���X���Rb�Έ�'}���2bPK�3�o/�-O�K�{1Ǘ��l�E�T�x4�6�;́I3��栳���L8�j:��q�8QkH'_�� 	ԉ�K�m�\$Œ�rD��O����g{9�e�pg�"
̓��4<�Q�N޲���&&0ly���rY�`��1B?�j����B�F�woB-�Ed���u�i#>�
Aj����3�SH����;nȚ%��J�2����-�$&�rH�.w{�FT`F��l��r�.�'x�O��6�(�J�N�%-]-e@؊@�,�����Q��9��?"��(��A֧���p� �>2�(;�%+�_.g"�﹔��7����L��>�A��C���V�{���2�ի@���[�L��Y��S�O��G|�p]�/��H[r:���M�"l�v�����`��N�%tb����p�D�Ls�#l�{�kV�&^i����n�E_L�i|�(�s��1�#N;�7�܆EN��s�-.'3k���o����� �i�dN�#>:��)bѡ���I�.�#�g�׉K���H��}xI�&� i�<9<�5M5E+"ˬ�]̝b���h�.�c�Ƽ��T�ef�:t����HĒ+��"\'�Z(������]�����F��KqMU�2�y��͊�����u	���`�罯��F7g}KK�։V1'�@�g�����Y�2��_�0D8�o\g��um��+>i�]��-Y�їw�K���Kyť.�F=��X�Owe��G\���FP<��x]yGBS�yt4�*h����] ��A�����1m8��W�O�y�$�Z����Ȳ ��q��	oXL���Al�����H�z�D���q;^T����X�z�C�"��a�a�}�\Zy���7��u8�9%����k���Ӷǯ�L ����3g���_;?*cA�8D�`�~�[��jE	��Z8d��da-��o��@������ C�����c�zR��^���0'W�t5��gf=�)n�]@Q���u(�P�[!à�=ձiH���M�V��J�r�6�ZS�x�آA����Cs����7�\�!�J��0���'��A�/\���T�F� �7j���1y\�� �86M����Kf&�W+F�\�f�gM 5��;%	]���Qmb-'�w@�.b�Hp�3��*/�,��I/�����@8�M����