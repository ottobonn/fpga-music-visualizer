library verilog;
use verilog.vl_types.all;
entity bel_fft_core is
    generic(
        word_width      : integer := 16;
        config_num      : integer := 1;
        stage_num       : integer := 4;
        twiddle_rom_max_awidth: integer := 8;
        fft_size        : integer := 256;
        fft_size1       : integer := 0;
        fft_size2       : integer := 0;
        fft_size3       : integer := 0;
        has_butterfly2  : integer := 1
    );
    port(
        clk_i           : in     vl_logic;
        rst_i           : in     vl_logic;
        butterfly_generic_adr_o: out    vl_logic_vector(31 downto 0);
        butterfly_generic_dat_re_i: in     vl_logic_vector;
        butterfly_generic_dat_re_o: out    vl_logic_vector;
        butterfly_generic_dat_im_i: in     vl_logic_vector;
        butterfly_generic_dat_im_o: out    vl_logic_vector;
        butterfly_generic_wr_o: out    vl_logic;
        butterfly_generic_rd_o: out    vl_logic;
        butterfly_generic_ack_i: in     vl_logic;
        butterfly_generic_err_i: in     vl_logic;
        butterfly2_adr_o: out    vl_logic_vector(31 downto 0);
        butterfly2_dat_re_i: in     vl_logic_vector;
        butterfly2_dat_re_o: out    vl_logic_vector;
        butterfly2_dat_im_i: in     vl_logic_vector;
        butterfly2_dat_im_o: out    vl_logic_vector;
        butterfly2_wr_o : out    vl_logic;
        butterfly2_rd_o : out    vl_logic;
        butterfly2_ack_i: in     vl_logic;
        butterfly2_err_i: in     vl_logic;
        butterfly4_adr_o: out    vl_logic_vector(31 downto 0);
        butterfly4_dat_re_i: in     vl_logic_vector;
        butterfly4_dat_re_o: out    vl_logic_vector;
        butterfly4_dat_im_i: in     vl_logic_vector;
        butterfly4_dat_im_o: out    vl_logic_vector;
        butterfly4_wr_o : out    vl_logic;
        butterfly4_rd_o : out    vl_logic;
        butterfly4_ack_i: in     vl_logic;
        butterfly4_err_i: in     vl_logic;
        copy_adr_o      : out    vl_logic_vector(31 downto 0);
        copy_dat_re_i   : in     vl_logic_vector;
        copy_dat_re_o   : out    vl_logic_vector;
        copy_dat_im_i   : in     vl_logic_vector;
        copy_dat_im_o   : out    vl_logic_vector;
        copy_wr_o       : out    vl_logic;
        copy_rd_o       : out    vl_logic;
        copy_ack_i      : in     vl_logic;
        copy_err_i      : in     vl_logic;
        ctrl_adr_i      : in     vl_logic_vector(9 downto 0);
        ctrl_dat_i      : in     vl_logic_vector(31 downto 0);
        ctrl_dat_o      : out    vl_logic_vector(31 downto 0);
        ctrl_bsel_i     : in     vl_logic_vector(3 downto 0);
        ctrl_wr_i       : in     vl_logic;
        ctrl_rd_i       : in     vl_logic;
        ctrl_ack_o      : out    vl_logic;
        ctrl_err_o      : out    vl_logic;
        tw_adr          : out    vl_logic_vector;
        tw_rd           : out    vl_logic;
        tw_re           : in     vl_logic_vector;
        tw_im           : in     vl_logic_vector;
        tw_cfg_sel      : out    vl_logic_vector;
        event_o         : out    vl_logic;
        int_o           : out    vl_logic;
        user_o          : out    vl_logic_vector(31 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of word_width : constant is 1;
    attribute mti_svvh_generic_type of config_num : constant is 1;
    attribute mti_svvh_generic_type of stage_num : constant is 1;
    attribute mti_svvh_generic_type of twiddle_rom_max_awidth : constant is 1;
    attribute mti_svvh_generic_type of fft_size : constant is 1;
    attribute mti_svvh_generic_type of fft_size1 : constant is 1;
    attribute mti_svvh_generic_type of fft_size2 : constant is 1;
    attribute mti_svvh_generic_type of fft_size3 : constant is 1;
    attribute mti_svvh_generic_type of has_butterfly2 : constant is 1;
end bel_fft_core;
